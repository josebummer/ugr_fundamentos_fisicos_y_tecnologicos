��  CCircuit��  CSerializeHack           ��  CPart            ���  CBattery��  CValue  ��    2V          @      �? V �� 	 CTerminal  �(�)        f�s��@�M��@�  �  �(	)        ���?�?�G���@?    ��4        ��      �� 	 CVoltRail
�  Kisw    2V(           @      �? V �  |p�q               @f��MbP?    tl|t         ����     ��  CEarth�  hxi�       	         &��Mbp�    [�s�         ��      ��  CCurrent
�  7Q__    4mA(    ����Mbp?      �?mA �  h8iM         X��C�@&��Mbp�  �  hdiy                &��Mbp?    `Lpd         ��      �� 	 CResistor
�  (H$    6k        p�@      �?k  �  D(Y)        X��C�@�G���@?  �  (-)        ���?�?�G���@�    ,$D,        ��      �
�  ��$    4k        @�@      �?k  �  �(�)     
  ���j�J$��3#�%�l�  �  x(�)        X��C�@�3#�%�l?    �$�,    "    ��      ��  C741��  COpampSupply�� 
 CDummyPart  �8�    (�  �8�      ��    14V            ,@      �? V       ,�      �? V % �   ��        f�s��@          �   ��        �3��@          �  ,�A�     
  ���j�J$��)&�%�l?    �,�     +      ��    ��  ��%       	         ����h?    �$�,     /    ��      �
�  ����    1k          @�@      �?k  �  ����         �3��@����h?  �  ���                ����h�    ����     2    ��      �
�  ����    3k        p�@      �?k  �  ����        �3��@����h�  �  ����       �3��'@����h?    ����    6    ��      �
�  Hh$    4k        @�@      �?k  �  d(y)        f�s��@�M��@?  �  8(M)        ��zA�j�?�M��@�    L$d,    :    ��      $�&�(�  0�P�    (�  0�P�      (�(�    14V            ,@      �? V       ,�      �? V < �  �-�       S����          �  �-�        ��zA�j�?          �  D�Y�       �3��'@����h�    ,�D�    @      ��    ��  ��%      	 	         f���MbP?    �$,     D    ��      �
�  ����    1mA(    ����MbP?      �?mA �  ���     	           f���MbP�  �  ����        S����f���MbP?    �� �    G    ��      �
�  ����    5k          ��@      �?k  �  ����         ��zA�j�?e���MbP?  �  ����       S����e���MbP�    ����     K    ��      �
�  �Z�h    1mA   ����MbP?      �?mA �  �p�q      	        @f��MbP�  �  �p�q        ��zA�j�?f��MbP?    �h�x    O    ��      �
�  ��$    2k        @�@      �?k  �  �(�)        ��zA�j�?�����X�  �  �(�)              @�����X?    �$�,    S    ��      �
�  +!S/    4V(          @      �? V �  \(q)              @�����X�    T$\,     W    ����                 ���  CWire  ()      Y�  �(�)      Y�  x(�)      Y�  ���      Y�  ��       Y�  �(9)      Y�  �(�q       Y�  ���      Y�  ����       Y�  �(�)      Y�  p(�)      Y�  �p��       Y�  �p�q      Y�  X���      Y�  ����       Y�  ����      Y�  ���      Y�  ���      Y�  ����       Y�  ����      Y�  �(��       Y�  h(y)      Y�  X(i)      Y�  h(i9       Y�  �(�)     
 Y�  �(��      
 Y�  @���     
             �                         [    Z   O     q       p  Z  " " r # o # ' ' + k + , j , - - t / 3 / 2 i 2 3 3 / 6 6 h 7 g 7 : : \ ; _ ; = = @ a @ A ^ A B B g D G D G G D H a H K e K L L b O  O P P f S S c T d T W W d   \  : n K ^ ] A c ; _ f b @ L H S ` W T ` ] P e B 7 6 i h j 2 , l + m k n l [ m p #  q o  " s r t - s            �$s�        @     +        @            @    "V  (      �8                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 