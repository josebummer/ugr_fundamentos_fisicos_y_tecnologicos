��  CCircuit��  CSerializeHack           ��  CPart              ���  CEarth�� 	 CTerminal  �X�m                 �&�Mb`�    �l�t         ��      �
�  � � %                             � $� ,         ��      �� 	 CResistor��  CValue  �n�|    3k        p�@      �?k  
�  ����       Kk�O�!�1K�3�  
�  p���     
         �!�1K�3?    �|��        ��      �� 	 CVoltRail�  Ks    6V(          @      �? V 
�  |�              @w�ȤYv�    t|         ����     ��  ��     2k        @�@      �?k  
�  	       ^�v8+N���]5Ar�  
�  ��	              @��]5Ar?    �        ��      ��  CCurrent�  �:�H    1mA   ����MbP?      �?mA 
�  �P	Q       ^�v8+N�WrMNbP�  
�  �P�Q              @WrMNbP?    �H�X        ��      ��  CBattery�  l� ��     9V         "@      �? V 
�  ��	     	   Q��c�X@�d���r�  
�  `u	       ^�v8+N���.�r?    t� �    $    ��      ��  �� �    3k        p�@      �?k  
�  �	       G��7,N��d���r�  
�  ��	     	   Q��c�X@�d���r?    ��    (    ��      ��  x>�L    6k        p�@      �?k  
�  �P�Q       G��7,N�D����J�  
�  hP}Q       ^�v8+N�D����J?    |L�T    ,    ��      ��  C741��  COpampSupply�� 
 CDummyPart  `l�z    2�  `���      X�X�    14V            ,@      �? V       ,�      �? V / 
�  H�]�       ^�v8+N�          
�  H�]�       Kk�O�          
�  t���       G��7,N���,�Yv?    \zt�     5      ��    ��  o	�    2mA(    ����Mb`?      �?mA 
�  ���        '�Z.��&�Mb`�  
�  ��1                �&�Mb`?    ��     :    ��      ��  ����    2k        @�@      �?k  
�  ���       Kk�O��1K�3?  
�  ����       '�Z.��1K�3�    ����    >    ��      ��  P�p�    1k        @�@      �?k  
�  l���       '�Z.���t��b?  
�  @�U�       �V[(O���t��b�    T�l�    B    ��      .�0�2�  � ��    2�  � ��      � �� �    8V             @      �? V        �      �? V D 
�  � �� �                          
�  � �� �     
         �          
�  � ��       �V[(O���t��b?    � �� �    H      ��    ��  c �� �    -2V(           �      �? V 
�  � �� �     
         �!�1K�3�    � �� �     M    ����                   ���  CWire  HPiQ      O�  8PIQ      O�  HPI�       O�  ��Q       O�  ��       O�  ��      O�  ��	      O�  P9Q      O�  89Q       O�  8a	      O�  9	      O�  ��	     	 O�   P	Q      O�  �PQ      O�   Q       O�  P	�       O�  ��	�      O�  � �� �     
 O�  � �� �      
 O�  � �q�     
 O�  (�I�      O�  (�)�       O�  (�)�       O�  ��)�      O�   �)�      O�  �A�      O�  �0�Y       O�  ����      O�  ����      O�  ����       O�  � ��        O�  � �� �      O�  � �� �      
               �                             j   n    g  c    U   Z  V    W   S   $ $ [ % Y % ( ( ^ ) [ ) , , ] - P - 1 1 5 R 5 6 d 6 7 7 ` : m : ; ; j > > h ? l ? B B k C i C E E H o H I p I J J i M M a Q - W R P 5 T   V U  S T   X Y Q Z %  X $ ) ] _ , ^ ( \ \ ` 7 _ M p c a b  f 6 g d e h  e > f J C ;  B m k ? l : o  n H b I            �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 