��  CCircuit��  CSerializeHack           ��  CPart              ���  C741��  COpampSupply�� 
 CDummyPart  0�P�    �  0P      (�(�    14V            ,@      �? V       ,�      �? V 	 �� 	 CTerminal   -     
   +�k  @          �  �-�        jJ���@          �  D�Y�       HT�n�'@ �D�J�    ,�D          ��    ��  CEarth�  (()=                        �    <3D         ��      ��  CBattery��  CValue  � �    8V(           @      �? V �  (�)�                @���Mb`�  �  ()!                ���Mb`?    �4         ��      ��  CCurrent�  ���    2mA(    ����Mb`?      �?mA �  ��!     
   +�k  @���Mb`�  �  ����         jJ���@���Mb`?    ���        ��      �� 	 CResistor�  ��$    2k        @�@      �?k  �  �(�)     
   +�k  @���Mb`?  �  p(�)                ���Mb`�    �$�,    $    ��      !��  ����    1k        @�@      �?k  �  ����        jJ���@���Mb`�  �  p���               @���Mb`?    ����    (    ��      ��  �P�e       	         ��D�J?    �dl     +    ��      !��  �)�7    5k          ��@      �?k  �  ��%         `ph>�@��D�J?  �  �<�Q                ��D�J�    �$�<     .    ��      ��  ����    3mA   �~j�t�h?      �?mA �  ����        ��{�@�ҡt�h�  �  ����       �@��a���ҡt�h?    ����    2    ��      �
��  h���    �  h���      `�`�    14V            ,@      �? V       ,�      �? V 4 �  P�e�        ��{�@          �  P�e�        `ph>�@          �  |���        ��|��? �3K�EM?    d�|�     8      ��    !��  ����    10k        ��@      �?k  �  ����        `ph>�@��D�J�  �  p���       HT�n�'@��D�J?    ����    =    ��      !��  P&p4    3k        p�@      �?k  �  l8�9        ��|��?�Y7K�EM�  �  @8U9        ��{�@�Y7K�EM?    T4l<    A    ��      !��  �&�4    4k        @�@      �?k  �  �8�9        ��{�@���Ba?  �  �8�9       �@��a�����Ba�    �4�<    E    ��      !��   &@4    0.50k        @@      �?k  �  <8Q9       �@��a���Y7K�EM�  �  8%9             ��Y7K�EM?    $4<<    I    ��      �� 	 CVoltRail�  �1�?    -4V(          �      �? V �  �8�9             ��Y7K�EM�    �4�<     N    ����                   ���  CWire  X�q�      P�   1      
 P�  �01     
 P�  ��       P�  ���      P�  ((q)      P�  (�q�      P�  (�)�       P�  ( ))       P�  � �1      
 P�  �0�1     
 P�  ����       P�  ����      P�  �(�1      
 P�  8�Q�      P�  8�9�       P�  ��9�      P�  ���       P�  ����      P�  �Q�      P�  ���      P�  �89      P�  h���      P�  h8i�       P�  P8i9      P�  h8�9      P�  ����      P�  �8��       P�  �8�9      P�  8�       P�  8A9      P�  �89                    �                               R   T    Q  V   X    Y   Z   \   $ $ ^ % V % ( ( ] ) W ) + / + . b . / / + 2 2 e 3 g 3 5 5 8 d 8 9 _ 9 : : k = = c > Q > A A m B o B E E f F j F I I i J p J N N p  >  S Z R U  \ T Y % X ) W     [ ^ S ]   ( U $ [ ` 9 _ a b ` c . = a n 8 2 d E n h 3 j g I h i F : l m k A l o e f B N J            �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 