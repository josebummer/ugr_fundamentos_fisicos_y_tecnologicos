��  CCircuit��  CSerializeHack           ��  CPart              ���  CCurrent��  CValue  /�W�    1mA(    ����MbP?      �?mA �� 	 CTerminal  `�a�                ��,�MbP�  �  `�a�       	 �_�J��@��,�MbP?    X�h�        ��      �� 	 CResistor
�  h� ��     3k        p�@      �?k  �  �� ��        !�&�$@�US�8a?  �  X� m�      
   y͘��@�US�8a�    l� ��         ��      �
�  �� ��     0.50k        @@      �?k  �  �� ��        !�&�$@ĪsB�?  �  x� ��       	 �1���?ĪsB��    �� ��         ��      ��  CBattery
�  D� l�     2V          @      �? V �  8� M�      
   y͘��@x��aB��  �  d� y�         �1���?ĪsB�?    L� d�         ��      �� 	 CVoltRail
�  I;W    4V(          @      �? V �  @8AM               @            <LDT         ����     ��  C741��  COpampSupply�� 
 CDummyPart  h�    %�  h/�=      ``    15V            .@      �? V       .�      �? V " �  Pe     
   y͘��@          �  P(e)              @          �  | �!       !�&�$@��r�_*��    d|/     (      ��    �
�  �� ��     1.5k        p�@      �?k  �  �� ��      
   y͘��@4Uq�zn{?  �  �� ��        ��o/�4Uq�zn{�    �� ��     -    ��      �
�  (    1k        @�@      �?k  �  $9     
   y͘��@�;�ρ��?  �  �       � L�
 ��;�ρ���    $    1    ��      �
�  �� ��     3k        p�@      �?k  �  �� ��        � L�
 ����c�E�  �  �� ��        ��o/����c�E?    �� ��     5    ��      �
�  L� t�     2V          @      �? V �  @� U�       	 ��o/�kG�t{p�  �  l� ��        ��o/��D��{p?    T� l�     9    ��      �
�  � 0�     2k        @�@      �?k  �  ,� A�        ��o/�kG�t{p?  �   � �        HJۛ�/(�kG�t{p�    � ,�     =    ��      �
�  @� `�     3k        p�@      �?k  �  \� q�        ��o/��&��O�`?  �  0� E�        HJۛ�/(��&��O�`�    D� \�     A    ��      !�#�%�  �� �
    %�  �'�5      ��    15V            .@      �? V       .�      �? V C �  ��       ��o/�          �  � �!       HJۛ�/�          �  ��       � L�
 �pD�c��?    �
�'     G      ��    ��  CEarth�  ����       	         Vt��h�    s���     L    ��      J��  8�9�      	 	         Vt��h�    +�C�     N    ��      �
�  [y{�    1k          @�@      �?k  �  �`�u       	 HJۛ�/�Vt��h�  �  ����                Vt��h?    |t��     Q    ��      �
�  y3�    2k          @�@      �?k  �  8`9u        HJۛ�/�Vt��h�  �  8�9�     	           Vt��h?    4t<�     U    ��      �
�  PNp\    1k        @�@      �?k  �  l`�a       HJۛ�/�Vt��h?  �  @`Ua       HJۛ�/�Vt��h�    T\ld    Y    ��      �
�  �N\    1k        @�@      �?k  �  `)a       HJۛ�/�Vt��x?  �  �`�a       HJۛ�/(�Vt��x�    �\d    ]    ��      J��  `�a�       	         ��,�MbP?    S�k�     `    ��      !�#�%�  �D�R    %�  �o�}      �X�X    15V            .@      �? V       .�      �? V a �  �X�Y        �����@          �  �h�i        �_�J��@          �  �`�a       HJۛ�/(�������?    �R�o     e      ��    �
�  ;a[o    4k          @�@      �?k  �  `Ha]       	 �����@��,�MbP?  �  `ta�        �_�J��@��,�MbP�    \\dt     j    ��      �
�  ;![/    5k          ��@      �?k  �  `a       	       (@��,�MbP?  �  `4aI        �����@��,�MbP�    \d4     n    ��      �
�  3� [�     12V(          (@      �? V �  `� a	             (@��,�MbP�    \� d�     r    ����                   ���  CWire  �� �!       t�  �� ��        t�  �� ��       t�  8� Y�      
 t�  8� 9�       
 t�  8� 9      
 t�  � �!      t�  @(Q)      t�  @(A9       t�  ��      t�  8Q     
 t�  �� 9�      
 t�  �� ��       t�  �� ��        t�  ��      t�  �� �       t�  �� ��       t�  �� ��       t�  p� ��       t�   � �        t�   � �        t�  �� �       t�  �� �a       t�  �`�a      t�  �`�a      t�   � 1�       t�  p� q       t�  p�      t�  0 �!      t�  0 1a       t�  (`1a      t�  0`9a      t�  8`Aa      t�  �h��       t�  `���      t�  �H�Y       t�  `H�I                    �                              `  k    w  x    v     y       }   $ $ (  ( ) | ) * * { - - � . � . 1 1 z 2 ~ 2 5 5 � 6 � 6 9 = 9 : : � = = 9 > � > A A � B � B D D G � G H � H I I � L R L N V N Q Y Q R R L U � U V V N Y Y Q Z � Z ] ] � ^ � ^ `  ` b b e � e f � f g g � j o j k k � n r n o o � r r n v {  w  u z  � x y  * u } ) |   � 2 1 ( -  : . � � I � � ~ 5 � � 6 � � � � > � � � � � g � � ^ � B A � � G � H � � ] � � U � Z f �  � � e j �            �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 