��  CCircuit��  CSerializeHack           ��  CPart              ���  CCurrent��  CValue  ��$�    2mA   ����Mb`?      �?mA �� 	 CTerminal  �1�       �^ۙ'@���Mb`�  �  ���        �dXE��ܿ���Mb`?    ��        ��      ��  CBattery
�  � Q� _    6V(          @      �? V �  8	M         �4����?Y+pMb`?  �  d	y       	�rX����L١Nb`�    � Ld         ��      ��  CEarth�  �`�u                             �t�|         ��      ��  C741��  COpampSupply�� 
 CDummyPart  �"    �  �?M      �(�(    14V            ,@      �? V       ,�      �? V  �  �(�)        �dXE��ܿ          �  �8�9                          �  �01       }�t��'@ Y~t�x�    �"�?           ��    �� 	 CResistor
�  S9sG    5k          ��@      �?k  �  x y5         �4����?Y+pMb`�  �  xLya       �^ۙ'@Y+pMb`?    t4|L     $    ��      !�
�  S�s�    4k          @�@      �?k  �  x�y�        �^ۙ'@��~�S��=  �  x�y	       }�t��'@��~�S���    t�|�     (    ��      !�
�  ���    2k        @�@      �?k  �  �!�       }�t��'@��;t�x?  �  ����        �dXE��ܿ��;t�x�    ���    ,    ��      !�
�  P�p�    1k        @�@      �?k  �  l���        �dXE��ܿUCxdMbp?  �  @�U�       	�rX���UCxdMbp�    T�l�    0    ��      �
�  � �� �    6mA(    �~j�t�x?      �?mA �  �	                ��d�t�x�  �  �	�        	�rX�����d�t�x?     ��    4    ��      ��  0	E                 ��d�t�x?    � DL     7    ��                    ���  CWire  ����       9�  ����      9�  0�y�      9�  x`y�       9�  x�y�       9�   y!      9�   	9       9�  x	�       9�  @0y1      9�  0A1      9�  @�A1       9�   �A�      9�  xy1       9�  �8�a       9�  �8�9      9�  �(�)      9�  ���)       9�  ����      9�  ����      9�  �A�      9�  �	�       9�  	1                     �                              <  ;   @    A  G     I   H      C $ ? $ % % = ( > ( ) ) F , , E - K - 0 0 L 1 M 1 4 4 O 5 N 5 7 O 7 L J :   > % < = ( @ $ ?   M C F   D E B , D ) B H  G  J  K I : - 0 ; N 1 A 5 4 7            �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 