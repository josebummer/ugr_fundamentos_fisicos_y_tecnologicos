��  CCircuit��  CSerializeHack           ��  CPart              ��� 	 CVoltRail��  CValue  ����    -7V         �      �? V �� 	 CTerminal  ����      	       �>�����%�    ����        ����     �� 	 CResistor
�  X�x�    1.2k        ��@      �?k  �  t���             �>�����%?  �  H�]�       ��H�X��>�����%�    \�t�        ��      �
�  �#�    0.40k           y@      �?k  �  (�)�        ��H�X���P/D�v?  �  (�)�       ǅ�f��"��P/D�v�    $�,�         ��      �
�  �#    0.20k           i@      �?k  �  (�)�       	 ǅ�f��"��P/D�v?  �  ()!       �$�[��$��P/D�v�    $�,         ��      �
�  ����    0.60k        ��@      �?k  �  ����       ��H�X���	O��u�  �  ����     	  �{�y���	O��u?    ����        ��      ��  C741��  COpampSupply�� 
 CDummyPart  `�    #�  `-�;      XX    15V            .@      �? V       .�      �? V   �  H(])       �$�[��$�          �  H]       ǅ�f��"�          �  t �!     
        *@            \t-    &      ��    ��  CCurrent
�  $�L�    1mA   ����MbP?      �?mA �  D�Y�       d�M���^}��MbP�  �  �-�        0M����^}��MbP?    ,�D�    ,    ��      �!�#�  ��    #�  �/�=      ��    15V            .@      �? V       .�      �? V . �  ��       d�M���          �  �(�)             �          �  � �!       �$�[��$��x/D�v?    ��/     2      ��    ��  CBattery
�  'D5    1V         �?      �? V �  @%A                ѥ��^��  �  <@QA             ��~�M�>    $4<L    8    ��      ��  CEarth�  � H� ]                 �?�|Ya`�    � \d     <    ��      �
�  Ss'    4k          @�@      �?k  �  x y        d�M����~�M�>  �  x,yA             ��~�M��    t|,     ?    ��      �
�  S�s�    3k          p�@      �?k  �  x�y�      	  �{�y��J=�^�aP�  �  x�y�       d�M���J=�^�aP?    t�|�     C    ��      �
�  � � '    1k          @�@      �?k  �  �  �          0M����`�j��a`�  �  � ,� A                `�j��a`?    � � ,     G    ��      �
�  � �� �    2k          @�@      �?k  �  � �� �      	 	 �{�y��d�3$�`P�  �  � �� �        0M����d�3$�`P?    � �� �     K    ��      �
�  � �� �    3k        p�@      �?k  �  � �� �     	  �{�y��=�{��Mk�  �  � �� �      	       @=�{��Mk?    � �� �    O    ��      �
�  s �� �    6V(          @      �? V �  � �� �              @=�{��Mk�    � �� �     S    ����                   ���  CWire  (�I�      U�  H�I       U�  (�I�      U�  ((I)      U�  ( ))       U�  � )!      U�  x���     	 U�  ����       U�  ��)�      U�  X�y�      U�  � ��      U�  � @� I       U�  � @A      U�  P@yA      U�  x@�A      U�  �(�A       U�  ���       U�  x���      U�  x�y�       U�  x�y       U�  � �y�     	 U�  � ��                      �                                   V   ^    X      [   ]  \  " " & Y & ' W ' ( (   , , _ - ` - / / 2 f 2 3 e 3 4 4 [ 8 b 8 9 9 c < a < ? i ? @ @ d C j C D D h G k G H H b K O K L L ` O O j P S P S S P   X '  W Z &  Y 4 Z C  ^  ] V , D k - H < a 8 9 @ c e 3 d g 2 i f _ g h ? K \ L G            �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 