��  CCircuit��  CSerializeHack           ��  CPart              ���  C741��  COpampSupply�� 
 CDummyPart  ����    �  ����      ����    14V            ,@      �? V       ,�      �? V 	 �� 	 CTerminal  ����        �H9���=          �  ����     	        (@          �  ����             (@            ����          ��    �� 	 CResistor��  CValue  �'    6k          p�@      �?k  �   	         �H9���= ���#�<  �  ,	A     
            ���#��    ,         ��      ��  CEarth�  h	}      
            ���#�<    �|�         ��      ��  8�X�    9k        ��@      �?k  �  T�i�        �H9���=          �  (�=�        �H9���=            <�T�        ��      �� 	 CVoltRail�  �AO    12V(          (@      �? V �  L	a     	        (@szj�t�h�    DL    #    ����     ��  �y�    4k          @�@      �?k  �  `	u      	 	       (@szj�t�h?  �  �	�        �H9���=szj�t�h�    t�     &    ��      ��  CCurrent�  ����    3mA   �~j�t�h?      �?mA �  ����        �<U4U?owj�t�h�  �  ����        �H9���=owj�t�h?    ����    +    ��      ��  (6HD    1k        @�@      �?k  �  DHYI        �<U4U?P`�Jbp�  �  H-I      	 9�7� @P`�Jbp?    ,DDL    /    ��      ��  CBattery�  �/=    2V          @      �? V �  �H�I        9�7� @R�tKbp?  �  HI        9�7� @P`�Jbp�    �<T    4    ��      1��  � �#�    1V(          �?      �? V �  0�1�              "@�v�!Pb`?  �  0�1�               @~�,�Mb`�    $�<�     8    ��       ��  � �� �    9V(          "@      �? V �  ��             "@�4w�s�x�    � ��     <    ����     (��  d2�@    3mA   �~j�t�h?      �?mA �  �H�I        9�7� @?���t�h�  �  XHmI       犣���?���t�h?    l@�P    ?    ��      �
��   � �    �   � �      ����    14V            ,@      �? V       ,�      �? V A �  ����        9�7� @          �  ����        [����@          �  �)�        �<U4U?c�@I�|?    ���     E      ��    ��  �h�}                 �Hh%NbP?    �|��     I    ��      (��  �)�7    1mA(    ����MbP?      �?mA �  �<�Q                �Hh%NbP�  �  ��%         [����@�Hh%NbP?    �$�<    L    ��      ��  h���    3k        p�@      �?k  �  ����        9�7� @Π�DbP�  �  X�m�             "@Π�DbP?    l���    P    ��      ��  h���    2k        @�@      �?k  �  � �        [����@ Ih%NbP�  �  X m               @ Ih%NbP?    l��    T    ��      ��  y+�    5k          ��@      �?k  �  0`1u        犣���?���t�h�  �  0�1�             "@?���t�h?    ,t4�     X    ��      ��  )+7    8k          @�@      �?k  �  01%                @����MbP?  �  0<1Q                ����MbP�    ,$4<     \    ��      ��  0p1�                 ����MbP?    #�;�     _    ��                    ���  CWire  ����       a�  ��	�      a�  �	       a�  �)�      a�  ��	�      a�  �	�       a�  h���      a�  ����     	 a�  �`��      	 a�  `�a     	 a�  @	i      
 a�  �H��       a�  �H��       a�  ����      a�  (���      a�  XH�I      a�  �H�I      a�   �1�      a�   �!�       a�  �!�      a�  0�1�       a�  0 Y      a�  0�1       a�  0�1�       a�  ����       a�  ����      a�  ����      a�  �H�I      a�  0HYI      a�  0H1a       a�  ����      a�  ���       a�  �P�i       a�  � �       a�  � �      a�  0�Y�      a�  0 1       a�  0P1q                     �                               h   i       d    l  l    h  e  # # k & # & ' ' g + o + , , f / / q 0 5 0 4 r 4 5 5 0 8 v 8 9 9 x < < u ? ? } @ ~ @ B B E | E F � F G G p I � I L L � M � M P P { Q � Q T T � U w U X  X Y Y y \ � \ ] ] � _ � _ , c b d c  f  b g ' e   j  k i & j   q o } { p + G m / m n 4 t Y s u < t � 8 � U 9 w s v n | P z z E ? r  @ ~ X � F � � L I � M T � y Q x \ ] _            �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 