��  CCircuit��  CSerializeHack           ��  CPart    H   H     ���  C741��  COpampSupply�� 
 CDummyPart  h���    �  h���      `�`�    15V            .@      �? V       .�      �? V 	 �� 	 CTerminal  P�e�        T����@          �  P�e�     	   �>4���@          �  |���             *@            d�|�          ��    �� 	 CResistor��  CValue  ���    3k          p�@      �?k  �  ��      	   �>4���@{�MbP?  �  ��        T����@{�MbP�    ��         ��      ��  ��    3k        p�@      �?k  �  ��        T����@{�MbP?  �  ��               @{�MbP�    ��        ��      ��  CEarth�  h�i�       	         C}t�h?    [�s�         ��      ��  CBattery�  3Y[g    2V(           @      �? V �  h@iU                @C}t�h?  �  hli�                C}t�h�    \Ttl     #    ��      ��  ��    2k        @�@      �?k  �  �	               @�?WMb`�  �  ��        �>4���@�?WMb`?    ��    '    ��      ��  @�`�    2k        @�@      �?k  �  \�q�     	   �>4���@ɃU�NbP�  �  0�E�             $@ɃU�NbP?    D�\�    +    ��      ��  @`    2k        @�@      �?k  �  \q        �>4���@▣NNb`�  �  0E             $@▣NNb`?    D\    /    ��       ��  k���    2V(           @      �? V �  ����      	   �>4���@  �{��>  �  ����        �>4���@�A<9{�>    ����     3    ��      �� 	 CVoltRail�  � �� �    10V(          $@      �? V �  � ��             $@�Xγu�h�    � �� �     8    ����         H   H     ���  CWire  ��      	 :�  ���     	 :�  �Q�     	 :�  ����      	 :�  p���     	 :�  P�Q�       :�  �Q�      :�  P�Q�      	 :�  �       :�  �      :�  h�      :�  hiA       :�  i      :�  ��      :�  ���       :�  p�      :�  �       :�  1      :�  ��       :�  �1�          H   H     �    H   H         H   H        @   B       =    C   D  E   $  # F # $ $  ' ' G ( H ( + + ? , N , / / J 0 L 0 3 > 3 4 4 I 8 8 M <  > ; ; B ? 3 + <  A  @ =  A D  C F  G # ' E I ( 4 J / H 8 L K 0 N K M ,  
          �$s�        @     +        @            @    "V  (      �h                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 